nameserver 172.24.170.29
nameserver 172.24.170.30
search india.ti.com
