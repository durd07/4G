domain india.ti.com broadcast
